// ============================================================================
// Tang Primer 25K 用 VGA トップモジュール
// ============================================================================
// ボード: Tang Primer 25K (Gowin GW5A-LV25MG121)
// 機能: 白黒VGA出力 (640x480@60Hz)
// クロック: 27MHz (オンボード) → そのままVGAに使用
// 出力: HSYNC, VSYNC, R, G, B (白黒なので全て同じ信号)
// ============================================================================

module VGA_BW_top(
    // クロックとリセット
    input  wire clk,            // 27MHz システムクロック (Tang Primer 25K オンボード)
    input  wire reset_btn,      // リセットボタン (Active High)
    
    // VGA出力
    output wire vga_hsync,      // VGA 水平同期信号
    output wire vga_vsync,      // VGA 垂直同期信号
    output wire vga_r,          // VGA 赤信号
    output wire vga_g,          // VGA 緑信号
    output wire vga_b           // VGA 青信号
);

    // ========================================================================
    // クロック設定
    // ========================================================================
    // Tang Primer 25Kは27MHzのオンボードクロックを搭載
    // VGA 640x480@60Hzの標準クロックは25.175MHz
    // 
    // 【オプション1】27MHzをそのまま使用 (簡易版・初心者向け)
    //   - 標準より約7%速いが、ほとんどのモニターで動作する
    //   - 設定不要で簡単
    //   - 現在のコードはこちらを使用
    //
    // 【オプション2】PLLで25.175MHzを生成 (正確・上級者向け)
    //   - Gowin IP Core GeneratorでPLLを生成
    //   - 下記のコメントアウト部分を有効化
    //   - より正確なVGAタイミングが得られる
    // ========================================================================
    
    wire clk_vga;
    
    // オプション1: 27MHzをそのまま使用 (デフォルト)
    assign clk_vga = clk;
    
    // オプション2: PLL使用 (使う場合は以下のコメントを外す)
    // Gowin_rPLL pll_inst (
    //     .clkout(clk_vga),       // 25.175MHz 出力
    //     .clkin(clk)             // 27MHz 入力
    // );

    // ========================================================================
    // VGA コアモジュール インスタンス化
    // ========================================================================
    
    wire video_signal;          // 白黒映像信号 (1=白, 0=黒)
    
    VGA_BW_simple vga_core (
        .clk_25mhz  (clk_vga),      // VGAクロック (27MHz)
        .reset      (reset_btn),    // リセット
        .hsync      (vga_hsync),    // 水平同期出力
        .vsync      (vga_vsync),    // 垂直同期出力
        .video      (video_signal)  // 映像信号出力
    );

    // ========================================================================
    // 白黒映像をRGB出力に接続
    // ========================================================================
    // 白黒(グレースケール)の場合、同じ信号をR/G/B全てに接続
    // video_signal = 1 のとき → R=G=B=1 → 白
    // video_signal = 0 のとき → R=G=B=0 → 黒
    
    assign vga_r = video_signal;
    assign vga_g = video_signal;
    assign vga_b = video_signal;

endmodule
