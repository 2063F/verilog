module question9
